module ArbTop(
    input                clk,
    
);






endmodule