module ArbTop(
    input                CLK,
    input                ASynReset_N,

);






endmodule